module plot

struct BarData {
	
}