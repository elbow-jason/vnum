module linalg

#flag -lopenblas -llapack
#include "cblas.h"
#include "lapacke.h"
