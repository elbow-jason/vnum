module la

#flag -framework Accelerate
#include "Accelerate/Accelerate.h"
