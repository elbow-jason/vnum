module vnum
