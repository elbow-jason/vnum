module vnum