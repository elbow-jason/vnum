module linalg

#flag -framework Accelerate
#include "Accelerate/Accelerate.h"
