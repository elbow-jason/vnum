module nn
