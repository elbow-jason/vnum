module fft

#flag -lfftw3
#include "fftw3.h"
