module vnum

pub const (
	VERSION = '0.1'
)