module plot
